module LightLED(
  input   clock,
  input   reset,
  output  io_led
);
  assign io_led = 1'h1; // @[LightLED.scala 18:12]
endmodule
